* Inverter for 23M1117 with 200 + 2 x 17 = 234ps delay.

*including model files for pMOS and nMOS

.include models-180nm.txt

*defining a parameter in order to scale the geometry of pMOS and nMOS

.param w_p=1.740 w_n=0.595
.param l_p=0.18 l_n=0.18

*defining a circuit component that can be called multiple times
*formula used for Area: AD=AS= Wx2Lmin and Perimeter: PD=PS= 2x(W+2Lmin)
.subckt inv supply Inp Out
MP1 Out Inp Supply Supply cmosp 
+ L={1u*{l_p}} W={{w_p}*1u} AD = {2*{w_p}*{l_p}*{1p}} AS = {2*{w_p}*{l_p}*{1p}} PD = {2*({w_p}+2*{l_p})*1u} PS = {2*({w_p}+2*{l_p})*1u}
MN1 Out Inp 0      0      cmosn
+ L={1u*{l_n}} W={{w_n}*1u} AD = {2*{w_n}*{l_n}*{1p}} AS = {2*{w_n}*{l_n}*{1p}} PD = {2*({w_n}+2*{l_n})*1u} PS = {2*({w_p}+2*{l_n})*1u}
.ends

* Main Supply
vdd supply 0 dc 1.8
*DUT
x1  supply Ck inv_out inv
* Load Capacitor
C1 inv_out 0 0.05pF
*DC Sweep from 0V to 1.8V with 0.1 steps of increments
Vck ck 0 1.8V
.DC VCk 0V 1.8V 1mV
.control
run
plot V(ck) V(inv_out)
*taking the derivative of the output curve to get to the slope of -1 in order to find noise margins
let dv = deriv(V(inv_out))

meas dc VIL find V(Ck) when dv=-1 fall=1
meas dc VIH find V(Ck) when dv=-1 rise=1
meas dc VOH find V(inv_out) when V(ck)=VIL  
meas dc VOL find V(inv_out) when V(ck)=VIH 

let highnoisemargin = VOH-VIH
print highnoisemargin
let lownoisemargin = VIL - VOL
print lownoisemargin

.endc
.end
