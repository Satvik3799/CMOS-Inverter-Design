* Inverter for 23M1117 with 200 + 2 x 17 = 234ps delay.

*including model files for pMOS and nMOS

.include models-180nm.txt

*defining a parameter in order to scale the geometry of pMOS and nMOS

.param w_p=1.740 w_n=0.595
.param l_p=0.18 l_n=0.18

*defining a circuit component that can be called multiple times
*formula used for Area: AD=AS= Wx2Lmin and Perimeter: PD=PS= 2x(W+2Lmin)
.subckt inv supply Inp Out
MP1 Out Inp Supply Supply cmosp 
+ L={1u*{l_p}} W={{w_p}*1u} AD = {2*{w_p}*{l_p}*{1p}} AS = {2*{w_p}*{l_p}*{1p}} PD = {2*({w_p}+2*{l_p})*1u} PS = {2*({w_p}+2*{l_p})*1u}
MN1 Out Inp 0      0      cmosn
+ L={1u*{l_n}} W={{w_n}*1u} AD = {2*{w_n}*{l_n}*{1p}} AS = {2*{w_n}*{l_n}*{1p}} PD = {2*({w_n}+2*{l_n})*1u} PS = {2*({w_p}+2*{l_n})*1u}
.ends

* Main Supply
vdd supply 0 dc 1.8
*DUT
x1  supply Ck inv_out inv
* Load Capacitor
C1 inv_out 0 0.05pF
*TRANSIENT ANALYSIS with pulse inputs
Vck  Ck   0 DC 0 PULSE(0 1.8 0nS 20pS 20pS 4nS 8.0nS)

* transient analysis with 1ps step size untill 35nS with 0nS of delay
.tran 1pS 35nS 0nS
.control
run
plot 4.0+V(Ck) V(inv_out)
meas tran inrise TRIG v(ck) VAL=0.18 RISE=2 TARG v(Ck) VAL=1.62 RISE=2
meas tran infall TRIG v(ck) VAL=1.62 FALL=2 TARG v(Ck) VAL=0.18 FALL=2
meas tran drise TRIG v(inv_out) VAL=0.18 RISE=2 TARG v(inv_out) VAL=1.62 RISE=2
meas tran dfall TRIG v(inv_out) VAL=1.62 FALL=2 TARG v(inv_out) VAL=0.18 FALL=2
.endc
.end
